// This module will mock the onboard CODEC for our FPGA
module codec(ADC_DAT, mclk, BCLK, DAC_DAT, I2C_SDAT, reset, SDI, SCLK, CH1, CH2, act);
  input DAC_DAT, mclk, reset, SDI, SCLK;
  output ADC_DAT, BCLK;
  //input signed 
  wire [0:32767] ADC_load;
  inout I2C_SDAT;
  output reg CH1, CH2;	//for testing purposes to determine if received byte is valid for address and sub-address
  output reg act;	// signals that the activate command has been received, allows reading/ writing of audio data
  // these registers are internal to the CODEC and represent the current
  // configuration
  reg[7:0] LLI, RLI, LHO, RHO, AAPC, DAPC, PDC, DAIF, SC, AC, RR; 
  
  reg state, nxt_state;
  reg[8:0] i2c_shift;
  reg[4:0] i2c_counter;
  reg SDI_old2, SDI_old, SCLK_old, SCLK_old2;
  reg[7:0] sub_addr;

  // audio storage wires and regs
  reg[32767:0] adc_data; // was 63:0
  reg[2047:0] dac_data;
  reg BCLK, ADC_DAT;
  reg[3:0] BCLK_counter;

  assign I2C_SDAT = ((i2c_counter == 5'h09) | (i2c_counter == 5'h12) | (i2c_counter == 5'h1b)) ? i2c_shift[0] : 1'bz; 
  // I2C_SDAT should be assigned conditionally to high when a byte is successfully received
  always@(posedge SCLK, negedge reset) begin
    if(!reset) begin
      state = 1'b0;
      SDI_old2 = 1'b1;
      SDI_old = 1'b1;
      SCLK_old = 1'b1;
      SCLK_old2 = 1'b1;
    end
    else begin
      state = nxt_state;
      SDI_old2 = SDI_old;
      SDI_old = SDI;
      SCLK_old2 = SCLK_old;
      SCLK_old = SCLK;
    end
  end

  always@(posedge SCLK, negedge reset) begin
    if(!reset) begin
      i2c_shift = 9'h1FF;
      i2c_counter = 5'h00;
      sub_addr = 8'h00;
      CH1 = 1'b0;
      CH2 = 1'b0;
      // set codec registers to default values from datasheet
      LLI = 8'h97;
      RLI = 8'h97;
      LHO = 8'h79;
      RHO = 8'h79;
      AAPC = 8'h0a;
      DAPC = 8'h08;
      PDC = 8'h9F;
      DAIF = 8'h0a;
      SC = 8'h00;
      AC = 8'h00;
      RR = 8'hFF;
      act = 1'b0;
    end
    else if((state == 1'b0)) begin
      i2c_counter = 5'h00;
      CH1 = 1'b0;
      CH2 = 1'b0;
    end
    else if(state == 1'b1) begin
      i2c_counter = i2c_counter + 1;
      i2c_shift = {i2c_shift[7:0], SDI};
      /*if((i2c_counter < 5'h08) | (i2c_counter > 5'h08 && i2c_counter < 5'h11) | (i2c_counter > 5'h11 && i2c_counter < 5'h1a)) begin
	      //i2c_counter = i2c_counter + 1;
	      nxt_state = 1'b1;
	      //i2c_shift = {i2c_shift[7:0], SDI};
      end*/
      if(i2c_counter == 5'h09) begin //ACK1
	//i2c_counter = i2c_counter + 1;
	//i2c_shift = {i2c_shift[7:0], SDI};
	//nxt_state = 1'b1;
	CH1 = (i2c_shift[8:1] == 8'h34) ? 1'b1 : 1'b0;

      end
      else if(i2c_counter == 5'h12) begin
      	//i2c_counter = i2c_counter + 1;
      	//i2c_shift = {i2c_shift[7:0], SDI};
      	//nxt_state = 1'b1;
      	sub_addr = i2c_shift[8:1];
      	CH2 = (i2c_shift[1] != 1'b1 && i2c_shift[8:1] <= 8'h14) ? 1'b1 : 1'b0; // checks for valid sub-address
      end
      else if(i2c_counter == 5'h1a) begin
	//i2c_counter = i2c_counter + 1;
	//i2c_shift = {i2c_shift[7:0], SDI};
	//nxt_state = 1'b1;
	// store data into codec register based on sub address, will not
	// store on an invalid address
	if(sub_addr == 8'h00) begin
	  LLI = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h02) begin
	  RLI = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h04) begin
	  LHO = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h06) begin
	  RHO = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h08) begin
	  AAPC = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h0a) begin
	  DAPC = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h0c) begin
	  PDC = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h0e) begin
	  DAIF = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h10) begin
	  SC = i2c_shift[7:0];
	end
	else if(sub_addr == 8'h12) begin
	  AC = i2c_shift[7:0];
	  act = 1'b1;
	end
	else if(sub_addr == 8'h14) begin
	  RR = i2c_shift[7:0];
	end
	      
      end
    end
  end

  always@(posedge SCLK, negedge reset, SDI) begin
    if(!reset) begin
      nxt_state = 1'b0;
      //i2c_shift = 9'h1FF;
      //i2c_counter = 5'h00;
      
    end
    else begin
      case(state)
	1'b0: begin
	  if(((SDI == 1'b0) && (SCLK == 1'b1) && (SDI_old2 == 1'b1))) begin //start bit
	    nxt_state = 1'b1;
	  end
	end
	1'b1: begin
	  if(((SDI == 1'b1) && (SCLK == 1'b1) && (SDI_old2 == 1'b0) && (i2c_counter >= 5'h1d))) begin //should only return to wait state once stop condition reached
	    nxt_state = 1'b0;
	    //i2c_counter = 5'h00;
	  end
	  /*else begin // only check these if posedge of SCLK
	    if((i2c_counter < 5'h08) | (i2c_counter > 5'h08 && i2c_counter < 5'h11) | (i2c_counter > 5'h11 && i2c_counter < 5'h1a)) begin
	      //i2c_counter = i2c_counter + 1;
	      nxt_state = 1'b1;
	      //i2c_shift = {i2c_shift[7:0], SDI};
	    end
	    else if(i2c_counter == 5'h08) begin //ACK1
	      //i2c_counter = i2c_counter + 1;
	      //i2c_shift = {i2c_shift[7:0], SDI};
	      nxt_state = 1'b1;
	      CH1 = (i2c_shift[8:1] == 8'h34) ? 1'b1 : 1'b0;

	    end
	    else if(i2c_counter == 5'h11) begin
	      //i2c_counter = i2c_counter + 1;
	      //i2c_shift = {i2c_shift[7:0], SDI};
	      nxt_state = 1'b1;
	      sub_addr = i2c_shift[8:1];
	      CH2 = (i2c_shift[1] != 1'b1 && i2c_shift[8:1] <= 8'h14) ? 1'b1 : 1'b0; // checks for valid sub-address
	    end
	    else if(i2c_counter == 5'h1a) begin
	      //i2c_counter = i2c_counter + 1;
	      //i2c_shift = {i2c_shift[7:0], SDI};
	      nxt_state = 1'b1;
	      // store data into codec register based on sub address, will not
	      // store on an invalid address
	      if(sub_addr == 8'h00) begin
		LLI = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h02) begin
		RLI = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h04) begin
		LHO = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h06) begin
		RHO = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h08) begin
		AAPC = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h0a) begin
		DAPC = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h0c) begin
		PDC = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h0e) begin
		DAIF = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h10) begin
		SC = i2c_shift[8:1];
	      end
	      else if(sub_addr == 8'h12) begin
		AC = i2c_shift[8:1];
		act = 1'b1;
	      end
	      else if(sub_addr == 8'h14) begin
		RR = i2c_shift[8:1];
	      end
	      
	    end
	    
  	  end*/
	  
	end
	default: begin
	  //nxt_state = 1'b0;
	  //CH1 = 1'b0;
	  //CH2 = 1'b0;
	end
      endcase
    end
  end

  // audio memory 
  always@(posedge mclk, negedge reset) begin
    if(!reset) begin
      BCLK_counter = 4'h0;
      BCLK = 1'b0;
    end
    else if(BCLK_counter == 4'he) begin
      BCLK_counter = 4'h0;
      BCLK = ~BCLK;
    end
    else begin
      BCLK_counter = BCLK_counter + 1;
    end
  end

  always@(posedge BCLK, negedge reset) begin
    if(!reset) begin
      adc_data = ADC_load;//64'h010147563d90143f;	//default starting audio data, loops on itself
      dac_data = 2048'd0;	//received data starts as empty
      ADC_DAT = 1'b0;
    end
    else if(act) begin
      ADC_DAT = adc_data[63];
      adc_data = {adc_data[32766:0], adc_data[32767]};
      dac_data = {dac_data[2046:0], DAC_DAT};
    end
  end

  assign ADC_load = 32768'b00000000000000000000000001101010000000001101010100000001001111000000000110100001000000100000001000000010010111110000001010110110000000110000011000000011010100000000001110010010000000111100110000000011111111010000010000100101000001000100010000000100010110010000010001100100000001000110010100000100010111000000010001001010000001000010111000000100000010010000001111011100000000111010011100000011011010010000001100100101000000101101101000000010100010100000001000110100000000011101101100000001100000000000000100100010000000001100010000000000011001100000000000000111111111111010110011111111010100111111111011111110111111101010110111111110011000101111111000011101111111011101111111111101101010011111110101111011111111010101010111111101001110011111110100100110111111010001110011111101000111001111110100100111111111010011101111111101010110001111110101111111111111011010111111111101111010001111111000101000111111100111000111111110110000001111111100010101111111110111000011111111110100000000000000110011000000001001100100000001000000100000000101101010000000011101001000000010001110110000001010100000000000110000001100000011011000110000001110111101000001000001001000000100011000000000010010101000000001001110011100000101000111100000010101001101000001010111001100000101100011110000010110100001000001011010101000000101101010000000010110011101000001011000100000000101011010010000010101000001000001010001000000000100110110010000010010011000000001000101000000000100000000100000001110101111000000110101011100000010111110100000001010011100000000100011101100000001110110010000000101110111000000010001011000000000101101110000000001011010000000000000000111111111101011011111111101011110111111110001011011111110110101001111111010011010111111100110100011111110001111111111111000011110111111100000100011111101111110101111110111110110111111011111110011111110000011001111111000100101111111100100100011111110011101001111111010101001111111101110010111111111001010101111111101110100111111111100011000000000000111000000000001110111000000001101011100000001001110000000000110011100000000100000000000000010011001000000001011001000000000110010100100000011100001110000001111100010000001000011100000000100100010000000010011010010000001010001010100000101010011110000010110000010000001011010110000000101110011010000010111100100000001011111001000000101111101100000010111110000000001011110000000000101110001100000010110100011000001010111011000000101010000000000010100000100000001001011111000000100011100100000010000011111000000111100011100000011011010100000001100001001000000101010011000000010001111110000000111011001000000010111001100000001000011000000000010101000000000000100011111111111111010011111111110010000111111110011110011111110111100001111111010101001111111100110101011111110001100111111111000000101111111011110000011111101110001011111110110110010111111011010101011111101101010111111110110110111111111011100101111111101111010011111111000010000111111100100000111111110011110001111111010111000111111101111111011111111010010111111111110011101111111111111001100000000010011100000000010101011000000010000101000000001011010100000000111001010000000100010100100000010100001010000001011100000000000110011011000000011100001110000001111010100000001000001100100000100010110000000010010001110000001001011110100000100111000110000010100000000000001010001001100000101000111010000010100011100000001010001001000000100111111100000010011100001000001001011100100000100100010010000010001001111000001000000111100000011110001010000001101110110000000110001111100000010110001000000001001100011000000011111111000000001100101110000000100101110000000001100010000000000010110101111111111110000111111111000100111111111001001001111111011000100111111100110100011111110000100011111110111000001111111010111011111111101001101101111110011111011111111001100101011111100101000101111110010000100111111000110111111111100011001001111110001100011111111000110110011111100011111011111110010011001111111001011111011111100111011001111110100100000111111010101111011111101101000101111110111101101111111100011110011111110100100011111111011101010111111110100010111111111101000100000000000000000000000000101111000000000101110110000000100010110000000010110111100000001110001000000001000010011000000100101111000000010101000100000001011100000000000110001010000000011010000100000001101100111000000111000001100000011100101000000001110011101000000111001110000000011100100010000001101111100000000110101111000000011001101100000001100000101000000101100101000000010100010010000001000111111000000011110111100000001100110000000000100111100000000001101110000000000011101110000000000010000111111111010011011111111001111001111111011010010111111100110100111111110000000101111110110011101111111010011110011111100111000011111110010001010111111000011101111111011111100011111101110110001111110110111011111111011010001111111101100011111111110110000001011111010111011101111101011100100111110101110001111111010111011011111101100000000111110110001110111111011010000111111101101110010111110111010100011111011111001111111110000101100111111000111100111111100110010101111110100100000111111010111101111111101110101111111111000110110111111101001011011111110111101101111111101010101111111111011001000000000000011010000000001100011000000001011010100000001000000100000000101001000000000011000100000000001101111110000000111110000000000100001011100000010001101010000001001001001000000100101010100000010010101100000001001001110000000100011101100000010001000000000000111111011000000011100110100000001100101100000000101010111000000010001000000000000110001000000000001110000000000000001011111111111101110011111111101011000111111101111010011111110100011011111111000100111111111011100000111111101010110101111110011110111111111001001011011111100001110011111101111100001111110111000111011111011010000101111101011111100111110101100000011111010100010101111101001011101111110100011101011111010001000001111101000010000111110100000101011111010000011101111101000011100111110100011001111111010010101001111101001111110111110101011000111111010111010111111101100101110111110110111100011111011110010001111110000011110111111000111100111111100110101111111110100111000111111011001110011111110000000001111111001100100111111101100100011111111001010011111111110001001111111111110010000000000001110100000000010001100000000001101011000000001000110110000000101010111000000011000110000000001101110000000000111011011000000011111010000000010000001000000001000001010000000100000011000000001111110000000000111100010000000011100000100000001100110000000000101100110000000010010110000000000111010100000000010100010000000000101001111111111111111111111111110100110111111110100100111111110111010101111111010001001111111100010011111111101110001011111110101100100111111010000011011111100101010011111110001010001111110111111111011111011101100001111101101101000111110110010011111111010111100001111101010111111111110101001011111111010011110001111101001100011111110100101100011111010010101101111101001011111111110100111000111111010100011011111101010110011111110101110001011111011000110011111101101011000111110111010000011111011111011101111110001000011111111001001110111111100111111011111110101100000111111011100010111111110001011101111111010010110111111101111111011111111011001111111111111001101000000000011000000000000100100000000000011101011000000010100000000000001100011110000000111011000000000100001100000000010010100010000001010000001000000101010100000000010110001010000001011011001000000101110010000000010111001000000001011011010000000101100011100000010101010110000001010000101000000100101011100000010001000010000000111100011000000011001111000000001010100110000000100000010000000001010110100000000010101001111111111111001111111111001101011111111001111001111111011011110111111101000000011111110001001011111110111001100111111010111011011111101001001101111110011011011111111001001011111111100010110011111110000100100111110111111011111111011110100101111101110110110111110111010010011111011100110111111101110011100111110111010011111111011101111001111101111011011111111000000001111111100001101001111110001101110111111001011000011111100111110101111110101001010111111011010000111111101111111101111111001011111111111101100010011111111001010111111111110010110000000000000000000000000011010100000000011010101000000010011110000000001101000010000001000000010000000100101111100000010101101100000001100000110000000110101000000000011100100100000001111001100000000111111110100000100001001010000010001000100000001000101100100000100011001000000010001100101000001000101110000000100010010100000010000101110000001000000100100000011110111000000001110100111000000110110100100000011001001010000001011011010000000101000101000000010001101000000000111011011000000011000000000000001001000100000000011000100000000000110011000000000000001111111111110101100111111110101001111111110111111101111111010101101111111100110001011111110000111011111110111011111111111011010100111111101011110111111110101010101111111010011100111111101001001101111110100011100111111010001110011111101001001111111110100111011111111010101100011111101011111111111110110101111111111011110100011111110001010001111111001110001111111101100000011111111000101011111111101110000111111111101000000000000001100110000000010011001000000010000001000000001011010100000000111010010000000100011101100000010101000000000001100000011000000110110001100000011101111010000010000010010000001000110000000000100101010000000010011100111000001010001111000000101010011010000010101110011000001011000111100000101101000010000010110101010000001011010100000000101100111010000010110001000000001010110100100000101010000010000010100010000000001001101100100000100100110000000010001010000000001000000001000000011101011110000001101010111000000101111101000000010100111000000001000111011000000011101100100000001011101110000000100010110000000001011011100000000010110100000000000000001111111111010110111111111010111101111111100010110111111101101010011111110100110101111111001101000111111100011111111111110000111101111111000001000111111011111101011111101111101101111110111111100111111100000110011111110001001011111111001001000111111100111010011111110101010011111111011100101111111110010101011111111011101001111111111000110000000000001110000000000011101110000000011010111000000010011100000000001100111000000001000000000000000100110010000000010110010000000001100101001000000111000011100000011111000100000010000111000000001001000100000000100110100100000010100010101000001010100111100000101100000100000010110101100000001011100110100000101111001000000010111110010000001011111011000000101111100000000010111100000000001011100011000000101101000110000010101110110000001010100000000000101000001000000010010111110000001000111001000000100000111110000001111000111000000110110101000000011000010010000001010100110000000100011111100000001110110010000000101110011000000010000110000000000101010000000000001000111111111111110100111111111100100001111111100111100111111101111000011111110101010011111111001101010111111100011001111111110000001011111110111100000111111011100010111111101101100101111110110101010111111011010101111111101101101111111110111001011111111011110100111111110000100001111111001000001111111100111100011111110101110001111111011111110111111110100101111111111100111011111111111110011000000000100111000000000101010110000000100001010000000010110101000000001110010100000001000101001000000101000010100000010111000000000001100110110000000111000011100000011110101000000010000011001000001000101100000000100100011100000010010111101000001001110001100000101000000000000010100010011000001010001110100000101000111000000010100010010000001001111111000000100111000010000010010111001000001001000100100000100010011110000010000001111000000111100010100000011011101100000001100011111000000101100010000000010011000110000000111111110000000011001011100000001001011100000000011000100000000000101101011111111111100001111111110001001111111110010010011111110110001001111111001101000111111100001000111111101110000011111110101110111111111010011011011111100111110111111110011001010111111001010001011111100100001001111110001101111111111000110010011111100011000111111110001101100111111000111110111111100100110011111110010111110111111001110110011111101001000001111110101011110111111011010001011111101111011011111111000111100111111101001000111111110111010101111111101000101111111111010001000000000000000000000000001011110000000001011101100000001000101100000000101101111000000011100010000000010000100110000001001011110000000101010001000000010111000000000001100010100000000110100001000000011011001110000001110000011000000111001010000000011100111010000001110011100000000111001000100000011011111000000001101011110000000110011011000000011000001010000001011001010000000101000100100000010001111110000000111101111000000011001100000000001001111000000000011011100000000000111011100000000000100001111111110100110111111110011110011111110110100101111111001101001111111100000001011111101100111011111110100111100111111001110000111111100100010101111110000111011111110111111000111111011101100011111101101110111111110110100011111111011000111111111101100000010111110101110111011111010111001001111101011100011111110101110110111111011000000001111101100011101111110110100001111111011011100101111101110101000111110111110011111111100001011001111110001111001111111001100101011111101001000001111110101111011111111011101011111111110001101101111111010010110111111101111011011111111010101011111111110110010000000000000110100000000011000110000000010110101000000010000001000000001010010000000000110001000000000011011111100000001111100000000001000010111000000100011010100000010010010010000001001010101000000100101011000000010010011100000001000111011000000100010000000000001111110110000000111001101000000011001011000000001010101110000000100010000000000001100010000000000011100000000000000010111111111111011100111111111010110001111111011110100111111101000110111111110001001111111110111000001111111010101101011111100111101111111110010010110111111000011100111111011111000011111101110001110111110110100001011111010111111001111101011000000111110101000101011111010010111011111101000111010111110100010000011111010000100001111101000001010111110100000111011111010000111001111101000110011111110100101010011111010011111101111101010110001111110101110101111111011001011101111101101111000111110111100100011111100000111101111110001111001111111001101011111111101001110001111110110011100111111100000000011111110011001001111111011001000111111110010100111111111100010011111111111100100000000000011101000000000100011000000000011010110000000010001101100000001010101110000000110001100000000011011100000000001110110110000000111110100000000100000010000000010000010100000001000000110000000011111100000000001111000100000000111000001000000011001100000000001011001100000000100101100000000001110101000000000101000100000000001010011111111111111111111111111101001101111111101001001111111101110101011111110100010011111111000100111111111011100010111111101011001001111110100000110111111001010100111111100010100011111101111111110111110111011000011111011011010001111101100100111111110101111000011111010101111111111101010010111111110100111100011111010011000111111101001011000111110100101011011111010010111111111101001110001111110101000110111111010101100111111101011100010111110110001100111111011010110001111101110100000111110111110111011111100010000111111110010011101111111001111110111111101011000001111110111000101111111100010111011111110100101101111111011111110111111110110011111111111110011010000000000110000000000001001000000000000111010110000000101000000000000011000111100000001110110000000001000011000000000100101000100000010100000010000001010101000000000101100010100000010110110010000001011100100000000101110010000000010110110100000001011000111000000101010101100000010100001010000001001010111000000100010000100000001111000110000000110011110000000010101001100000001000000100000000010101101000000000101010011111111111110011111111110011010111111110011110011111110110111101111111010000000111111100010010111111101110011001111110101110110111111010010011011111100110110111111110010010111111111000101100111111100001001001111101111110111111110111101001011111011101101101111101110100100111110111001101111111011100111001111101110100111111110111011110011111011110110111111110000000011111111000011010011111100011011101111110010110000111111001111101011111101010010101111110110100001111111011111111011111110010111111111111011000100111111110010101111111111100101100000000000000000000000000110101000000000110101010000000100111100000000011010000100000010000000100000001001011111000000101011011000000011000001100000001101010000000000111001001000000011110011000000001111111101000001000010010100000100010001000000010001011001000001000110010000000100011001010000010001011100000001000100101000000100001011100000010000001001000000111101110000000011101001110000001101101001000000110010010100000010110110100000001010001010000000100011010000000001110110110000000110000000000000010010001000000000110001000000000001100110000000000000011111111111101011001111111101010011111111101111111011111110101011011111111001100010111111100001110111111101110111111111110110101001111111010111101111111101010101011111110100111001111111010010011011111101000111001111110100011100111111010010011111111101001110111111110101011000111111010111111111111101101011111111110111101000111111100010100011111110011100011111111011000000111111110001010111111111011100001111111111010000000000000011001100000000100110010000000100000010000000010110101000000001110100100000001000111011000000101010000000000011000000110000001101100011000000111011110100000100000100100000010001100000000001001010100000000100111001110000010100011110000001010100110100000101011100110000010110001111000001011010000100000101101010100000010110101000000001011001110100000101100010000000010101101001000001010100000100000101000100000000010011011001000001001001100000000100010100000000010000000010000000111010111100000011010101110000001011111010000000101001110000000010001110110000000111011001000000010111011100000001000101100000000010110111000000000101101000000000000000011111111110101101111111110101111011111111000101101111111011010100111111101001101011111110011010001111111000111111111111100001111011111110000010001111110111111010111111011111011011111101111111001111111000001100111111100010010111111110010010001111111001110100111111101010100111111110111001011111111100101010111111110111010011111111110001100000000000011100000000000111011100000000110101110000000100111000000000011001110000000010000000000000001001100100000000101100100000000011001010010000001110000111000000111110001000000100001110000000010010001000000001001101001000000101000101010000010101001111000001011000001000000101101011000000010111001101000001011110010000000101111100100000010111110110000001011111000000000101111000000000010111000110000001011010001100000101011101100000010101000000000001010000010000000100101111100000010001110010000001000001111100000011110001110000001101101010000000110000100100000010101001100000001000111111000000011101100100000001011100110000000100001100000000001010100000000000010001111111111111101001111111111001000011111111001111001111111011110000111111101010100111111110011010101111111000110011111111100000010111111101111000001111110111000101111111011011001011111101101010101111110110101011111111011011011111111101110010111111110111101001111111100001000011111110010000011111111001111000111111101011100011111110111111101111111101001011111111111001110111111111111100110000000001001110000000001010101100000001000010100000000101101010000000011100101000000010001010010000001010000101000000101110000000000011001101100000001110000111000000111101010000000100000110010000010001011000000001001000111000000100101111010000010011100011000001010000000000000101000100110000010100011101000001010001110000000101000100100000010011111110000001001110000100000100101110010000010010001001000001000100111100000100000011110000001111000101000000110111011000000011000111110000001011000100000000100110001100000001111111100000000110010111000000010010111000000000110001000000000001011010111111111111000011111111100010011111111100100100111111101100010011111110011010001111111000010001111111011100000111111101011101111111110100110110111111001111101111111100110010101111110010100010111111001000010011111100011011111111110001100100111111000110001111111100011011001111110001111101111111001001100111111100101111101111110011101100111111010010000011111101010111101111110110100010111111011110110111111110001111001111111010010001111111101110101011111111010001011111111110100010000000000000000000000000010111100000000010111011000000010001011000000001011011110000000111000100000000100001001100000010010111100000001010100010000000101110000000000011000101000000001101000010000000110110011100000011100000110000001110010100000000111001110100000011100111000000001110010001000000110111110000000011010111100000001100110110000000110000010100000010110010100000001010001001000000100011111100000001111011110000000110011000000000010011110000000000110111000000000001110111000000000001000011111111101001101111111100111100111111101101001011111110011010011111111000000010111111011001110111111101001111001111110011100001111111001000101011111100001110111111101111110001111110111011000111111011011101111111101101000111111110110001111111111011000000101111101011101110111110101110010011111010111000111111101011101101111110110000000011111011000111011111101101000011111110110111001011111011101010001111101111100111111111000010110011111100011110011111110011001010111111010010000011111101011110111111110111010111111111100011011011111110100101101111111011110110111111110101010111111111101100100000000000001101000000000110001100000000101101010000000100000010000000010100100000000001100010000000000110111111000000011111000000000010000101110000001000110101000000100100100100000010010101010000001001010110000000100100111000000010001110110000001000100000000000011111101100000001110011010000000110010110000000010101011100000001000100000000000011000100000000000111000000000000000101111111111110111001111111110101100011111110111101001111111010001101111111100010011111111101110000011111110101011010111111001111011111111100100101101111110000111001111110111110000111111011100011101111101101000010111110101111110011111010110000001111101010001010111110100101110111111010001110101111101000100000111110100001000011111010000010101111101000001110111110100001110011111010001100111111101001010100111110100111111011111010101100011111101011101011111110110010111011111011011110001111101111001000111111000001111011111100011110011111110011010111111111010011100011111101100111001111111000000000111111100110010011111110110010001111111100101001111111111000100111111111111001000000000000111010000000001000110000000000110101100000000100011011000000010101011100000001100011000000000110111000000000011101101100000001111101000000001000000100000000100000101000000010000001100000000111111000000000011110001000000001110000010000000110011000000000010110011000000001001011000000000011101010000000001010001000000000010100111111111111111111111111111010011011111111010010011111111011101010111111101000100111111110001001111111110111000101111111010110010011111101000001101111110010101001111111000101000111111011111111101111101110110000111110110110100011111011001001111111101011110000111110101011111111111010100101111111101001111000111110100110001111111010010110001111101001010110111110100101111111111010011100011111101010001101111110101011001111111010111000101111101100011001111110110101100011111011101000001111101111101110111111000100001111111100100111011111110011111101111111010110000011111101110001011111111000101110111111101001011011111110111111101111111101100111111111111100110100000000001100000000000010010000000000001110101100000001010000000000000110001111000000011101100000000010000110000000001001010001000000101000000100000010101010000000001011000101000000101101100100000010111001000000001011100100000000101101101000000010110001110000001010101011000000101000010100000010010101110000001000100001000000011110001100000001100111100000000101010011000000010000001000000000101011010000000001010100111111111111100111111111100110101111111100111100111111101101111011111110100000001111111000100101111111011100110011111101011101101111110100100110111111001101101111111100100101111111110001011001111111000010010011111011111101111111101111010010111110111011011011111011101001001111101110011011111110111001110011111011101001111111101110111100111110111101101111111100000000111111110000110100111111000110111011111100101100001111110011111010111111010100101011111101101000011111110111111110111111100101111111111110110001001111111100101011111111111001011000000000000000000000000001101010000000001101010100000001001111000000000110100001000000100000001000000010010111110000001010110110000000110000011000000011010100000000001110010010000000111100110000000011111111010000010000100101000001000100010000000100010110010000010001100100000001000110010100000100010111000000010001001010000001000010111000000100000010010000001111011100000000111010011100000011011010010000001100100101000000101101101000000010100010100000001000110100000000011101101100000001100000000000000100100010000000001100010000000000011001100000000000000111111111111010110011111111010100111111111011111110111111101010110111111110011000101111111000011101111111011101111111111101101010011111110101111011111111010101010111111101001110011111110100100110111111010001110011111101000111001111110100100111111111010011101111111101010110001111110101111111111111011010111111111101111010001111111000101000111111100111000111111110110000001111111100010101111111110111000011111111110100000000000000110011000000001001100100000001000000100000000101101010000000011101001000000010001110110000001010100000000000110000001100000011011000110000001110111101000001000001001000000100011000000000010010101000000001001110011100000101000111100000010101001101000001010111001100000101100011110000010110100001000001011010101000000101101010000000010110011101000001011000100000000101011010010000010101000001000001010001000000000100110110010000010010011000000001000101000000000100000000100000001110101111000000110101011100000010111110100000001010011100000000100011101100000001110110010000000101110111000000010001011000000000101101110000000001011010000000000000000111111111101011011111111101011110111111110001011011111110110101001111111010011010111111100110100011111110001111111111111000011110111111100000100011111101111110101111110111110110111111011111110011111110000011001111111000100101111111100100100011111110011101001111111010101001111111101110010111111111001010101111111101110100111111111100011000000000000111000000000001110111000000001101011100000001001110000000000110011100000000100000000000000010011001000000001011001000000000110010100100000011100001110000001111100010000001000011100000000100100010000000010011010010000001010001010100000101010011110000010110000010000001011010110000000101110011010000010111100100000001011111001000000101111101100000010111110000000001011110000000000101110001100000010110100011000001010111011000000101010000000000010100000100000001001011111000000100011100100000010000011111000000111100011100000011011010100000001100001001000000101010011000000010001111110000000111011001000000010111001100000001000011000000000010101000000000000100011111111111111010011111111110010000111111110011110011111110111100001111111010101001111111100110101011111110001100111111111000000101111111011110000011111101110001011111110110110010111111011010101011111101101010111111110110110111111111011100101111111101111010011111111000010000111111100100000111111110011110001111111010111000111111101111111011111111010010111111111110011101111111111111001100000000010011100000000010101011000000010000101000000001011010100000000111001010000000100010100100000010100001010000001011100000000000110011011000000011100001110000001111010100000001000001100100000100010110000000010010001110000001001011110100000100111000110000010100000000000001010001001100000101000111010000010100011100000001010001001000000100111111100000010011100001000001001011100100000100100010010000010001001111000001000000111100000011110001010000001101110110000000110001111100000010110001000000001001100011000000011111111000000001100101110000000100101110000000001100010000000000010110101111111111110000111111111000100111111111001001001111111011000100111111100110100011111110000100011111110111000001111111010111011111111101001101101111110011111011111111001100101011111100101000101111110010000100111111000110111111111100011001001111110001100011111111000110110011111100011111011111110010011001111111001011111011111100111011001111110100100000111111010101111011111101101000101111110111101101111111100011110011111110100100011111111011101010111111110100010111111111101000100000000000000000000000000101111000000000101110110000000100010110000000010110111100000001110001000000001000010011000000100101111000000010101000100000001011100000000000110001010000000011010000100000001101100111000000111000001100000011100101000000001110011101000000111001110000000011100100010000001101111100000000110101111000000011001101100000001100000101000000101100101000000010100010010000001000111111000000011110111100000001100110000000000100111100000000001101110000000000011101110000000000010000111111111010011011111111001111001111111011010010111111100110100111111110000000101111110110011101111111010011110011111100111000011111110010001010111111000011101111111011111100011111101110110001111110110111011111111011010001111111101100011111111110110000001011111010111011101111101011100100111110101110001111111010111011011111101100000000111110110001110111111011010000111111101101110010111110111010100011111011111001111111110000101100111111000111100111111100110010101111110100100000111111010111101111111101110101111111111000110110111111101001011011111110111101101111111101010101111111111011001000000000000011010000000001100011000000001011010100000001000000100000000101001000000000011000100000000001101111110000000111110000000000100001011100000010001101010000001001001001000000100101010100000010010101100000001001001110000000100011101100000010001000000000000111111011000000011100110100000001100101100000000101010111000000010001000000000000110001000000000001110000000000000001011111111111101110011111111101011000111111101111010011111110100011011111111000100111111111011100000111111101010110101111110011110111111111001001011011111100001110011111101111100001111110111000111011111011010000101111101011111100111110101100000011111010100010101111101001011101111110100011101011111010001000001111101000010000111110100000101011111010000011101111101000011100111110100011001111111010010101001111101001111110111110101011000111111010111010111111101100101110111110110111100011111011110010001111110000011110111111000111100111111100110101111111110100111000111111011001110011111110000000001111111001100100111111101100100011111111001010011111111110001001111111111110010000000000001110100000000010001100000000001101011000000001000110110000000101010111000000011000110000000001101110000000000111011011000000011111010000000010000001000000001000001010000000100000011000000001111110000000000111100010000000011100000100000001100110000000000101100110000000010010110000000000111010100000000010100010000000000101001111111111111111111111111110100110111111110100100111111110111010101111111010001001111111100010011111111101110001011111110101100100111111010000011011111100101010011111110001010001111110111111111011111011101100001111101101101000111110110010011111111010111100001111101010111111111110101001011111111010011110001111101001100011111110100101100011111010010101101111101001011111111110100111000111111010100011011111101010110011111110101110001011111011000110011111101101011000111110111010000011111011111011101111110001000011111111001001110111111100111111011111110101100000111111011100010111111110001011101111111010010110111111101111111011111111011001111111111111001101000000000011000000000000100100000000000011101011000000010100000000000001100011110000000111011000000000100001100000000010010100010000001010000001000000101010100000000010110001010000001011011001000000101110010000000010111001000000001011011010000000101100011100000010101010110000001010000101000000100101011100000010001000010000000111100011000000011001111000000001010100110000000100000010000000001010110100000000010101001111111111111001111111111001101011111111001111001111111011011110111111101000000011111110001001011111110111001100111111010111011011111101001001101111110011011011111111001001011111111100010110011111110000100100111110111111011111111011110100101111101110110110111110111010010011111011100110111111101110011100111110111010011111111011101111001111101111011011111111000000001111111100001101001111110001101110111111001011000011111100111110101111110101001010111111011010000111111101111111101111111001011111111111101100010011111111001010111111111110010110;



endmodule
